module igmv(OUT, ADDR, DATA1, DATA2_0, DATA2_1, DATA2_2, DATA2_3, DATA2_4, DATA2_5, DATA2_6, DATA2_7, DATA2_8, DATA2_9, Read, RD, ST, CLK, RST);
	output [319:0] OUT;
	output [3:0] ADDR;
	input [31:0] DATA1;
	input [31:0] DATA2_0;
	input [31:0] DATA2_1;
	input [31:0] DATA2_2;
	input [31:0] DATA2_3;
	input [31:0] DATA2_4;
	input [31:0] DATA2_5;
	input [31:0] DATA2_6;
	input [31:0] DATA2_7;
	input [31:0] DATA2_8;
	input [31:0] DATA2_9;
	output Read;
	output RD;
	input ST;
	input CLK;
	input RST;

	wire RD0;
	wire RD1;
	wire RD2;
	wire RD3;
	wire RD4;
	wire RD5;
	wire RD6;
	wire RD7;
	wire RD8;
	wire RD9;
	wire Read0;
	wire Read1;
	wire Read2;
	wire Read3;
	wire Read4;
	wire Read5;
	wire Read6;
	wire Read7;
	wire Read8;
	wire Read9;

	assign RD = RD0 & RD1 & RD2 & RD3 & RD4 & RD5 & RD6 & RD7 & RD8 & RD9 ;
	assign Read = Read0 & Read1 & Read2 & Read3 & Read4 & Read5 & Read6 & Read7 & Read8 & Read9 ;
	rowmult rowmult0(OUT[31:0], ST, RD0, CLK, RST, DATA1, DATA2_0, ADDR, Read0);
	defparam rowmult0.matrix_width = 11;
	defparam rowmult0.data_width = 32;
	defparam rowmult0.address_width = 4;
	rowmult rowmult1(OUT[63:32], ST, RD1, CLK, RST, DATA1, DATA2_1, ADDR, Read1);
	defparam rowmult1.matrix_width = 11;
	defparam rowmult1.data_width = 32;
	defparam rowmult1.address_width = 4;
	rowmult rowmult2(OUT[95:64], ST, RD2, CLK, RST, DATA1, DATA2_2, ADDR, Read2);
	defparam rowmult2.matrix_width = 11;
	defparam rowmult2.data_width = 32;
	defparam rowmult2.address_width = 4;
	rowmult rowmult3(OUT[127:96], ST, RD3, CLK, RST, DATA1, DATA2_3, ADDR, Read3);
	defparam rowmult3.matrix_width = 11;
	defparam rowmult3.data_width = 32;
	defparam rowmult3.address_width = 4;
	rowmult rowmult4(OUT[159:128], ST, RD4, CLK, RST, DATA1, DATA2_4, ADDR, Read4);
	defparam rowmult4.matrix_width = 11;
	defparam rowmult4.data_width = 32;
	defparam rowmult4.address_width = 4;
	rowmult rowmult5(OUT[191:160], ST, RD5, CLK, RST, DATA1, DATA2_5, ADDR, Read5);
	defparam rowmult5.matrix_width = 11;
	defparam rowmult5.data_width = 32;
	defparam rowmult5.address_width = 4;
	rowmult rowmult6(OUT[223:192], ST, RD6, CLK, RST, DATA1, DATA2_6, ADDR, Read6);
	defparam rowmult6.matrix_width = 11;
	defparam rowmult6.data_width = 32;
	defparam rowmult6.address_width = 4;
	rowmult rowmult7(OUT[255:224], ST, RD7, CLK, RST, DATA1, DATA2_7, ADDR, Read7);
	defparam rowmult7.matrix_width = 11;
	defparam rowmult7.data_width = 32;
	defparam rowmult7.address_width = 4;
	rowmult rowmult8(OUT[287:256], ST, RD8, CLK, RST, DATA1, DATA2_8, ADDR, Read8);
	defparam rowmult8.matrix_width = 11;
	defparam rowmult8.data_width = 32;
	defparam rowmult8.address_width = 4;
	rowmult rowmult9(OUT[319:288], ST, RD9, CLK, RST, DATA1, DATA2_9, ADDR, Read9);
	defparam rowmult9.matrix_width = 11;
	defparam rowmult9.data_width = 32;
	defparam rowmult9.address_width = 4;
endmodule

module igmv_tb();
	wire [31:0] DATA1;
	wire [31:0] DATA2_0;
	wire [31:0] DATA2_1;
	wire [31:0] DATA2_2;
	wire [31:0] DATA2_3;
	wire [31:0] DATA2_4;
	wire [31:0] DATA2_5;
	wire [31:0] DATA2_6;
	wire [31:0] DATA2_7;
	wire [31:0] DATA2_8;
	wire [31:0] DATA2_9;
	wire [3:0] ADDR;
	wire RD;
	wire [319:0] OUT;
	reg rST;
	reg rCLK;
	reg rRST;
	wire ST;
	wire CLK;
	wire RST;
	syncmemory mem0(.OUT_DATA(DATA2_0), .ADDR(ADDR), .RD(Read), .CLK(CLK), .RST(RST));
	defparam mem0.data_width = 32;
	defparam mem0.depth = 10;
	defparam mem0.address_width = 4;
	defparam mem0.input_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_0.bin";
	defparam mem0.output_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_0o.bin";
	syncmemory mem1(.OUT_DATA(DATA2_1), .ADDR(ADDR), .RD(Read), .CLK(CLK), .RST(RST));
	defparam mem1.data_width = 32;
	defparam mem1.depth = 10;
	defparam mem1.address_width = 4;
	defparam mem1.input_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_1.bin";
	defparam mem1.output_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_1o.bin";
	syncmemory mem2(.OUT_DATA(DATA2_2), .ADDR(ADDR), .RD(Read), .CLK(CLK), .RST(RST));
	defparam mem2.data_width = 32;
	defparam mem2.depth = 10;
	defparam mem2.address_width = 4;
	defparam mem2.input_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_2.bin";
	defparam mem2.output_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_2o.bin";
	syncmemory mem3(.OUT_DATA(DATA2_3), .ADDR(ADDR), .RD(Read), .CLK(CLK), .RST(RST));
	defparam mem3.data_width = 32;
	defparam mem3.depth = 10;
	defparam mem3.address_width = 4;
	defparam mem3.input_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_3.bin";
	defparam mem3.output_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_3o.bin";
	syncmemory mem4(.OUT_DATA(DATA2_4), .ADDR(ADDR), .RD(Read), .CLK(CLK), .RST(RST));
	defparam mem4.data_width = 32;
	defparam mem4.depth = 10;
	defparam mem4.address_width = 4;
	defparam mem4.input_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_4.bin";
	defparam mem4.output_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_4o.bin";
	syncmemory mem5(.OUT_DATA(DATA2_5), .ADDR(ADDR), .RD(Read), .CLK(CLK), .RST(RST));
	defparam mem5.data_width = 32;
	defparam mem5.depth = 10;
	defparam mem5.address_width = 4;
	defparam mem5.input_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_5.bin";
	defparam mem5.output_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_5o.bin";
	syncmemory mem6(.OUT_DATA(DATA2_6), .ADDR(ADDR), .RD(Read), .CLK(CLK), .RST(RST));
	defparam mem6.data_width = 32;
	defparam mem6.depth = 10;
	defparam mem6.address_width = 4;
	defparam mem6.input_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_6.bin";
	defparam mem6.output_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_6o.bin";
	syncmemory mem7(.OUT_DATA(DATA2_7), .ADDR(ADDR), .RD(Read), .CLK(CLK), .RST(RST));
	defparam mem7.data_width = 32;
	defparam mem7.depth = 10;
	defparam mem7.address_width = 4;
	defparam mem7.input_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_7.bin";
	defparam mem7.output_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_7o.bin";
	syncmemory mem8(.OUT_DATA(DATA2_8), .ADDR(ADDR), .RD(Read), .CLK(CLK), .RST(RST));
	defparam mem8.data_width = 32;
	defparam mem8.depth = 10;
	defparam mem8.address_width = 4;
	defparam mem8.input_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_8.bin";
	defparam mem8.output_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_8o.bin";
	syncmemory mem9(.OUT_DATA(DATA2_9), .ADDR(ADDR), .RD(Read), .CLK(CLK), .RST(RST));
	defparam mem9.data_width = 32;
	defparam mem9.depth = 10;
	defparam mem9.address_width = 4;
	defparam mem9.input_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_9.bin";
	defparam mem9.output_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_9o.bin";
	syncmemory mem_vector(.OUT_DATA(DATA1), .ADDR(ADDR), .RD(Read), .CLK(CLK), .RST(RST));
	defparam mem_vector.data_width = 32;
	defparam mem_vector.depth = 10;
	defparam mem_vector.address_width = 4;
	defparam mem_vector.input_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_vector.bin";
	defparam mem_vector.output_file = "d:/Work/dissertation_microprocessor/altera_projects/fpga_igmv/matrices/test_vectoro.bin";
	assign RST = rRST;
	assign CLK = rCLK;
	assign ST = rST;
igmv igmv1(OUT, ADDR, DATA1, DATA2_0, DATA2_1, DATA2_2, DATA2_3, DATA2_4, DATA2_5, DATA2_6, DATA2_7, DATA2_8, DATA2_9, Read, RD, ST, CLK, RST);
	always begin
		#5 rCLK = ~rCLK;
	end
	initial begin
		rCLK = 0;
		rST = 0;
		rRST = 0;
		#5 rRST = 1;
		#5 rRST = 0;
		#5 rST = 1;
		#5 rST = 0;
	end
endmodule
