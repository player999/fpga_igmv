library verilog;
use verilog.vl_types.all;
entity igmv_tb is
end igmv_tb;
